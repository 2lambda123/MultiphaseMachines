
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.MATH_REAL.all;
use ieee.std_logic_unsigned.all;


package array14bit_pkg is
  type array14bit is array (natural range <>) of std_logic_vector(13 downto 0);
end package;

package body array14bit_pkg is
end package body;

